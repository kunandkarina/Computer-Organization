module Shifter( result, leftRight, shamt, sftSrc  );
    
  output wire[31:0] result;

  input wire leftRight;
  input wire[4:0] shamt;
  input wire[31:0] sftSrc ;
  
  /*your code here*/ 
  wire [31:0] ls;
  wire [31:0] rs;
  
  and(rs[31], sftSrc[31], ~leftRight);
  and(rs[30], sftSrc[30], ~leftRight);
  and(rs[29], sftSrc[29], ~leftRight);
  and(rs[28], sftSrc[28], ~leftRight);
  and(rs[27], sftSrc[27], ~leftRight);
  and(rs[26], sftSrc[26], ~leftRight);
  and(rs[25], sftSrc[25], ~leftRight);
  and(rs[24], sftSrc[24], ~leftRight);
  and(rs[23], sftSrc[23], ~leftRight);
  and(rs[22], sftSrc[22], ~leftRight);
  and(rs[21], sftSrc[21], ~leftRight);
  and(rs[20], sftSrc[20], ~leftRight);
  and(rs[19], sftSrc[19], ~leftRight);
  and(rs[18], sftSrc[18], ~leftRight);
  and(rs[17], sftSrc[17], ~leftRight);
  and(rs[16], sftSrc[16], ~leftRight);
  and(rs[15], sftSrc[15], ~leftRight);
  and(rs[14], sftSrc[14], ~leftRight);
  and(rs[13], sftSrc[13], ~leftRight);
  and(rs[12], sftSrc[12], ~leftRight);
  and(rs[11], sftSrc[11], ~leftRight);
  and(rs[10], sftSrc[10], ~leftRight);
  and(rs[9], sftSrc[9], ~leftRight);
  and(rs[8], sftSrc[8], ~leftRight);
  and(rs[7], sftSrc[7], ~leftRight);
  and(rs[6], sftSrc[6], ~leftRight);
  and(rs[5], sftSrc[5], ~leftRight);
  and(rs[4], sftSrc[4], ~leftRight);
  and(rs[3], sftSrc[3], ~leftRight);
  and(rs[2], sftSrc[2], ~leftRight);
  and(rs[1], sftSrc[1], ~leftRight);
  
  and(ls[31], sftSrc[30], leftRight);
  and(ls[30], sftSrc[29], leftRight);
  and(ls[29], sftSrc[28], leftRight);
  and(ls[28], sftSrc[27], leftRight);
  and(ls[27], sftSrc[26], leftRight);
  and(ls[26], sftSrc[25], leftRight);
  and(ls[25], sftSrc[24], leftRight);
  and(ls[24], sftSrc[23], leftRight);
  and(ls[23], sftSrc[22], leftRight);
  and(ls[22], sftSrc[21], leftRight);
  and(ls[21], sftSrc[20], leftRight);
  and(ls[20], sftSrc[19], leftRight);
  and(ls[19], sftSrc[18], leftRight);
  and(ls[18], sftSrc[17], leftRight);
  and(ls[17], sftSrc[16], leftRight);
  and(ls[16], sftSrc[15], leftRight);
  and(ls[15], sftSrc[14], leftRight);
  and(ls[14], sftSrc[13], leftRight);
  and(ls[13], sftSrc[12], leftRight);
  and(ls[12], sftSrc[11], leftRight);
  and(ls[11], sftSrc[10], leftRight);
  and(ls[10], sftSrc[9], leftRight);
  and(ls[9], sftSrc[8], leftRight);
  and(ls[8], sftSrc[7], leftRight);
  and(ls[7], sftSrc[6], leftRight);
  and(ls[6], sftSrc[5], leftRight);
  and(ls[5], sftSrc[4], leftRight);
  and(ls[4], sftSrc[3], leftRight);
  and(ls[3], sftSrc[2], leftRight);
  and(ls[2], sftSrc[1], leftRight);
  and(ls[1], sftSrc[0], leftRight);
  
  or(result[31], 0, ls[31]);
  or(result[30], rs[31], ls[30]);
  or(result[29], rs[30], ls[29]);
  or(result[28], rs[29], ls[28]);
  or(result[27], rs[28], ls[27]);
  or(result[26], rs[27], ls[26]);
  or(result[25], rs[26], ls[25]);
  or(result[24], rs[25], ls[24]);
  or(result[23], rs[24], ls[23]);
  or(result[22], rs[23], ls[22]);
  or(result[21], rs[22], ls[21]);
  or(result[20], rs[21], ls[20]);
  or(result[19], rs[20], ls[19]);
  or(result[18], rs[19], ls[18]);
  or(result[17], rs[18], ls[17]);
  or(result[16], rs[17], ls[16]);
  or(result[15], rs[16], ls[15]);
  or(result[14], rs[15], ls[14]);
  or(result[13], rs[14], ls[13]);
  or(result[12], rs[13], ls[12]);
  or(result[11], rs[12], ls[11]);
  or(result[10], rs[11], ls[10]);
  or(result[9], rs[10], ls[9]);
  or(result[8], rs[9], ls[8]);
  or(result[7], rs[8], ls[7]);
  or(result[6], rs[7], ls[6]);
  or(result[5], rs[6], ls[5]);
  or(result[4], rs[5], ls[4]);
  or(result[3], rs[4], ls[3]);
  or(result[2], rs[3], ls[2]);
  or(result[1], rs[2], ls[1]);
  or(result[0], rs[1], 0);
	
endmodule